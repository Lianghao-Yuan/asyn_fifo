package fifo_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import fifo_agent_pkg::*;
  `include "fifo_read_seq.svh"
  `include "fifo_write_seq.svh"
  `include "fifo_test.svh"

endpackage: fifo_test_pkg
